module Auto_LevelUp(
    iState_flag,
    iRST_level_ctrl,
    iLevel,

    orst
);